module fsmboothmult(
	input start,
	input valid,
	output prodload,
	output multload,
	output 
);




endmodule