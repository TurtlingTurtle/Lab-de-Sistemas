module boothmult(
	input[5:0] A,
	input[5:0] B,
	output[11:0] R
);

endmodule